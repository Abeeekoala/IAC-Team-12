module ALU #(
    DATA_WIDTH = 32
) (
    input logic     ALUop1,
    input logic     ALUop2,
    input logic     ALUctrl,
    output logic    ALUout,
    output logic    eq

);
    
endmodule