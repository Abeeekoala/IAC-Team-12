module top(
    input   logic           clk,
    input   logic           rst,
    output  logic           a0         
);



    
endmodule